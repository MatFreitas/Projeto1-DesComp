library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

--		  tmp(0)  := "0100000000001"; -- LDI 1
--        tmp(1)  := "0101100000000"; -- STA 0
--		  tmp(2)  := "0010100000000"; -- SOMA 0
--        tmp(3)  := "0101100000001"; -- STA 1
--		  tmp(4)  := "0001100000000"; -- LDA 0
--        tmp(5)  := "0101100000001"; -- STA 257
--        tmp(6)  := "0101100000010"; -- STA 258
--        tmp(7)  := "0100001010101"; -- LDI 85
--        tmp(8)  := "0101100000000"; -- STA 256
--        tmp(9)  := "0100010101010"; -- LDI 170
--        tmp(10) := "0101100000000"; -- STA 256 
--        tmp(11) := "0110000001011"; -- JMP 11
--        tmp(12) := "0000000000000";
--        tmp(13) := "0000000000000";
--        tmp(14) := "0000000000000";
--        tmp(15) := "0000000000000";
		  
		  
--		  tmp(0)  := "0001101000000"; -- LDA 320
--        tmp(1)  := "0101100100000"; -- STA 288
--		  tmp(2)  := "0001101000001"; -- LDA 321
--        tmp(3)  := "0101100100001"; -- STA 289
--		  tmp(4)  := "0001101000010"; -- LDA 322
--        tmp(5)  := "0101100100010"; -- STA 290
--        tmp(6)  := "0001101100000"; -- LDA 352
--        tmp(7)  := "0101100100101"; -- STA 293
--        tmp(8)  := "0001101100001"; -- LDA 353
--        tmp(9)  := "0101100100110"; -- STA 294
--        tmp(10) := "0001101100010"; -- LDA 354	
--        tmp(11) := "0101100100110"; -- STA 294
--        tmp(12) := "0001101100011"; -- LDA 355	
--        tmp(13) := "0101100000001"; -- STA 257	
--        tmp(14) := "0001101100100"; -- LDA 356	
--        tmp(15) := "0101100000010"; -- STA 258
--		  tmp(16) := "0110000000000"; -- JMP 0
		  
--		  tmp(0)  := "0100000000001"; -- LDI 1
--        tmp(1)  := "0101000000000"; -- STA 0
--		  tmp(2)  := "0010" & '0' & "0000" & "0000"; -- SOMA 0
--        tmp(3)  := "0101100100000"; -- STA 288
--		  tmp(4)  := "0010000000000"; -- SOMA 0
--        tmp(5)  := "0101100100001"; -- STA 289
--        tmp(6)  := "0010000000000"; -- SOMA 0	
--        tmp(7)  := "0101100100010"; -- STA 290	
--        tmp(8)  := "0010000000000"; -- SOMA 0	
--        tmp(9)  := "0101100100011"; -- STA 291	
--        tmp(10) := "0010000000000"; -- SOMA 0		
--        tmp(11) := "0101100100100"; -- STA 292	
--        tmp(12) := "0010000000000"; -- SOMA 0	
--        tmp(13) := "0101100100101"; -- STA 293		
--        tmp(14) := "0110000000010"; -- JMP 2		
--        tmp(15) := "0000000000000"; 
--		  tmp(16) := "0000000000000"; 

--		  tmp(0)  := "0001101000000"; -- LDA 320
--        tmp(1)  := "0101100100000"; -- STA 288
--		  tmp(2)  := "0001101000001"; -- LDA 321
--        tmp(3)  := "0101100100001"; -- STA 289
--		  tmp(4)  := "0001101000010"; -- LDA 322
--        tmp(5)  := "0101100100010"; -- STA 290			
--        tmp(6)  := "0001101100000"; -- LDA 352		
--        tmp(7)  := "0101100100011"; -- STA 291	
--        tmp(8)  := "0001101100001"; -- LDA 353	
--        tmp(9)  := "0101100100100"; -- STA 292		
--        tmp(10) := "0001101100010"; -- LDA 354		
--        tmp(11) := "0101100100101"; -- STA 293	
--        tmp(12) := "0001101100011"; -- LDA 355	
--        tmp(13) := "0101100000001"; -- STA 257	
--        tmp(14) := "0001101100100"; -- LDA 356		
--        tmp(15) := "0101100000010"; -- STA 258
--		  tmp(16) := "0110000000000"; -- JMP 0	
		  
		  tmp(0)  := "0100000000000"; -- LDI 0	
        tmp(1)  := "0101000000000"; -- STA 0	
		  tmp(2)  := "0101000000010"; -- STA 2	
        tmp(3)  := "0100000000001"; -- LDI 1	
		  tmp(4)  := "0101000000001"; -- STA 1	
        tmp(5)  := "0000000000000"; -- NOP			
        tmp(6)  := "0001101100000"; -- LDA 352		
        tmp(7)  := "1000000000000"; -- CEQ 0		
        tmp(8)  := "0111000001010"; -- JEQ 10	
        tmp(9)  := "1001000100000"; -- JSR 32		
        tmp(10) := "0000000000000"; -- NOP		
        tmp(11) := "0110000000101"; -- JMP 5	
        tmp(32) := "0101111111111"; -- STA 511	
        tmp(33) := "0001000000010"; -- LDA 2	
        tmp(34) := "0010000000001"; -- SOMA 1		
        tmp(35) := "0101000000010"; -- STA 2	
		  tmp(36) := "0101100000010"; -- STA 258	
		  tmp(37) := "1010000000000"; -- STA 258	
		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;